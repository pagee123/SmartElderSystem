module rx(
    input rx_pin,
    output  tx_pin
    );
 assign	tx_pin=rx_pin;
				
endmodule